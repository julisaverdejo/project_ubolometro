// Author: Julisa Verdejo Palacios
// Name: rom_volts.v
//
// Description: 


module rom_volts (
  input      [8:0] addr_i,
  output reg [11:0] rom_o
);

  always@(addr_i)  
    case(addr_i)
        0 : rom_o = 12'b000000000000; //0.000000
        1 : rom_o = 12'b000000000000; //0.000000
        2 : rom_o = 12'b000000000000; //0.000000
        3 : rom_o = 12'b000000000000; //0.000000
        4 : rom_o = 12'b000000000000; //0.000000
        5 : rom_o = 12'b000000000000; //0.000000
        6 : rom_o = 12'b000000000000; //0.000000
        7 : rom_o = 12'b000000000000; //0.000000
        8 : rom_o = 12'b000000000000; //0.000000
        9 : rom_o = 12'b000000000000; //0.000000
       10 : rom_o = 12'b000001111100; //0.100000
       11 : rom_o = 12'b000001111100; //0.100000
       12 : rom_o = 12'b000001111100; //0.100000
       13 : rom_o = 12'b000001111100; //0.100000
       14 : rom_o = 12'b000001111100; //0.100000
       15 : rom_o = 12'b000001111100; //0.100000
       16 : rom_o = 12'b000001111100; //0.100000
       17 : rom_o = 12'b000001111100; //0.100000
       18 : rom_o = 12'b000001111100; //0.100000
       19 : rom_o = 12'b000001111100; //0.100000
       20 : rom_o = 12'b000011111000; //0.200000
       21 : rom_o = 12'b000011111000; //0.200000
       22 : rom_o = 12'b000011111000; //0.200000
       23 : rom_o = 12'b000011111000; //0.200000
       24 : rom_o = 12'b000011111000; //0.200000
       25 : rom_o = 12'b000011111000; //0.200000
       26 : rom_o = 12'b000011111000; //0.200000
       27 : rom_o = 12'b000011111000; //0.200000
       28 : rom_o = 12'b000011111000; //0.200000
       29 : rom_o = 12'b000011111000; //0.200000
       30 : rom_o = 12'b000101110100; //0.300000
       31 : rom_o = 12'b000101110100; //0.300000
       32 : rom_o = 12'b000101110100; //0.300000
       33 : rom_o = 12'b000101110100; //0.300000
       34 : rom_o = 12'b000101110100; //0.300000
       35 : rom_o = 12'b000101110100; //0.300000
       36 : rom_o = 12'b000101110100; //0.300000
       37 : rom_o = 12'b000101110100; //0.300000
       38 : rom_o = 12'b000101110100; //0.300000
       39 : rom_o = 12'b000101110100; //0.300000
       40 : rom_o = 12'b000111110000; //0.400000
       41 : rom_o = 12'b000111110000; //0.400000
       42 : rom_o = 12'b000111110000; //0.400000
       43 : rom_o = 12'b000111110000; //0.400000
       44 : rom_o = 12'b000111110000; //0.400000
       45 : rom_o = 12'b000111110000; //0.400000
       46 : rom_o = 12'b000111110000; //0.400000
       47 : rom_o = 12'b000111110000; //0.400000
       48 : rom_o = 12'b000111110000; //0.400000
       49 : rom_o = 12'b000111110000; //0.400000
       50 : rom_o = 12'b001001101100; //0.500000
       51 : rom_o = 12'b001001101100; //0.500000
       52 : rom_o = 12'b001001101100; //0.500000
       53 : rom_o = 12'b001001101100; //0.500000
       54 : rom_o = 12'b001001101100; //0.500000
       55 : rom_o = 12'b001001101100; //0.500000
       56 : rom_o = 12'b001001101100; //0.500000
       57 : rom_o = 12'b001001101100; //0.500000
       58 : rom_o = 12'b001001101100; //0.500000
       59 : rom_o = 12'b001001101100; //0.500000
       60 : rom_o = 12'b001011101000; //0.600000
       61 : rom_o = 12'b001011101000; //0.600000
       62 : rom_o = 12'b001011101000; //0.600000
       63 : rom_o = 12'b001011101000; //0.600000
       64 : rom_o = 12'b001011101000; //0.600000
       65 : rom_o = 12'b001011101000; //0.600000
       66 : rom_o = 12'b001011101000; //0.600000
       67 : rom_o = 12'b001011101000; //0.600000
       68 : rom_o = 12'b001011101000; //0.600000
       69 : rom_o = 12'b001011101000; //0.600000
       70 : rom_o = 12'b001101100100; //0.700000
       71 : rom_o = 12'b001101100100; //0.700000
       72 : rom_o = 12'b001101100100; //0.700000
       73 : rom_o = 12'b001101100100; //0.700000
       74 : rom_o = 12'b001101100100; //0.700000
       75 : rom_o = 12'b001101100100; //0.700000
       76 : rom_o = 12'b001101100100; //0.700000
       77 : rom_o = 12'b001101100100; //0.700000
       78 : rom_o = 12'b001101100100; //0.700000
       79 : rom_o = 12'b001101100100; //0.700000
       80 : rom_o = 12'b001111100000; //0.800000
       81 : rom_o = 12'b001111100000; //0.800000
       82 : rom_o = 12'b001111100000; //0.800000
       83 : rom_o = 12'b001111100000; //0.800000
       84 : rom_o = 12'b001111100000; //0.800000
       85 : rom_o = 12'b001111100000; //0.800000
       86 : rom_o = 12'b001111100000; //0.800000
       87 : rom_o = 12'b001111100000; //0.800000
       88 : rom_o = 12'b001111100000; //0.800000
       89 : rom_o = 12'b001111100000; //0.800000
       90 : rom_o = 12'b010001011100; //0.900000
       91 : rom_o = 12'b010001011100; //0.900000
       92 : rom_o = 12'b010001011100; //0.900000
       93 : rom_o = 12'b010001011100; //0.900000
       94 : rom_o = 12'b010001011100; //0.900000
       95 : rom_o = 12'b010001011100; //0.900000
       96 : rom_o = 12'b010001011100; //0.900000
       97 : rom_o = 12'b010001011100; //0.900000
       98 : rom_o = 12'b010001011100; //0.900000
       99 : rom_o = 12'b010001011100; //0.900000
      100 : rom_o = 12'b010011011000; //1.000000
      101 : rom_o = 12'b010011011000; //1.000000
      102 : rom_o = 12'b010011011000; //1.000000
      103 : rom_o = 12'b010011011000; //1.000000
      104 : rom_o = 12'b010011011000; //1.000000
      105 : rom_o = 12'b010011011000; //1.000000
      106 : rom_o = 12'b010011011000; //1.000000
      107 : rom_o = 12'b010011011000; //1.000000
      108 : rom_o = 12'b010011011000; //1.000000
      109 : rom_o = 12'b010011011000; //1.000000
      110 : rom_o = 12'b010101010100; //1.100000
      111 : rom_o = 12'b010101010100; //1.100000
      112 : rom_o = 12'b010101010100; //1.100000
      113 : rom_o = 12'b010101010100; //1.100000
      114 : rom_o = 12'b010101010100; //1.100000
      115 : rom_o = 12'b010101010100; //1.100000
      116 : rom_o = 12'b010101010100; //1.100000
      117 : rom_o = 12'b010101010100; //1.100000
      118 : rom_o = 12'b010101010100; //1.100000
      119 : rom_o = 12'b010101010100; //1.100000
      120 : rom_o = 12'b010111010000; //1.200000
      121 : rom_o = 12'b010111010000; //1.200000
      122 : rom_o = 12'b010111010000; //1.200000
      123 : rom_o = 12'b010111010000; //1.200000
      124 : rom_o = 12'b010111010000; //1.200000
      125 : rom_o = 12'b010111010000; //1.200000
      126 : rom_o = 12'b010111010000; //1.200000
      127 : rom_o = 12'b010111010000; //1.200000
      128 : rom_o = 12'b010111010000; //1.200000
      129 : rom_o = 12'b010111010000; //1.200000
      130 : rom_o = 12'b011001001100; //1.300000
      131 : rom_o = 12'b011001001100; //1.300000
      132 : rom_o = 12'b011001001100; //1.300000
      133 : rom_o = 12'b011001001100; //1.300000
      134 : rom_o = 12'b011001001100; //1.300000
      135 : rom_o = 12'b011001001100; //1.300000
      136 : rom_o = 12'b011001001100; //1.300000
      137 : rom_o = 12'b011001001100; //1.300000
      138 : rom_o = 12'b011001001100; //1.300000
      139 : rom_o = 12'b011001001100; //1.300000
      140 : rom_o = 12'b011011001000; //1.400000
      141 : rom_o = 12'b011011001000; //1.400000
      142 : rom_o = 12'b011011001000; //1.400000
      143 : rom_o = 12'b011011001000; //1.400000
      144 : rom_o = 12'b011011001000; //1.400000
      145 : rom_o = 12'b011011001000; //1.400000
      146 : rom_o = 12'b011011001000; //1.400000
      147 : rom_o = 12'b011011001000; //1.400000
      148 : rom_o = 12'b011011001000; //1.400000
      149 : rom_o = 12'b011011001000; //1.400000
      150 : rom_o = 12'b011101000100; //1.500000
      151 : rom_o = 12'b011101000100; //1.500000
      152 : rom_o = 12'b011101000100; //1.500000
      153 : rom_o = 12'b011101000100; //1.500000
      154 : rom_o = 12'b011101000100; //1.500000
      155 : rom_o = 12'b011101000100; //1.500000
      156 : rom_o = 12'b011101000100; //1.500000
      157 : rom_o = 12'b011101000100; //1.500000
      158 : rom_o = 12'b011101000100; //1.500000
      159 : rom_o = 12'b011101000100; //1.500000
      160 : rom_o = 12'b011111000000; //1.600000
      161 : rom_o = 12'b011111000000; //1.600000
      162 : rom_o = 12'b011111000000; //1.600000
      163 : rom_o = 12'b011111000000; //1.600000
      164 : rom_o = 12'b011111000000; //1.600000
      165 : rom_o = 12'b011111000000; //1.600000
      166 : rom_o = 12'b011111000000; //1.600000
      167 : rom_o = 12'b011111000000; //1.600000
      168 : rom_o = 12'b011111000000; //1.600000
      169 : rom_o = 12'b011111000000; //1.600000
      170 : rom_o = 12'b100000111100; //1.700000
      171 : rom_o = 12'b100000111100; //1.700000
      172 : rom_o = 12'b100000111100; //1.700000
      173 : rom_o = 12'b100000111100; //1.700000
      174 : rom_o = 12'b100000111100; //1.700000
      175 : rom_o = 12'b100000111100; //1.700000
      176 : rom_o = 12'b100000111100; //1.700000
      177 : rom_o = 12'b100000111100; //1.700000
      178 : rom_o = 12'b100000111100; //1.700000
      179 : rom_o = 12'b100000111100; //1.700000
      180 : rom_o = 12'b100010111000; //1.800000
      181 : rom_o = 12'b100010111000; //1.800000
      182 : rom_o = 12'b100010111000; //1.800000
      183 : rom_o = 12'b100010111000; //1.800000
      184 : rom_o = 12'b100010111000; //1.800000
      185 : rom_o = 12'b100010111000; //1.800000
      186 : rom_o = 12'b100010111000; //1.800000
      187 : rom_o = 12'b100010111000; //1.800000
      188 : rom_o = 12'b100010111000; //1.800000
      189 : rom_o = 12'b100010111000; //1.800000
      190 : rom_o = 12'b100100110100; //1.900000
      191 : rom_o = 12'b100100110100; //1.900000
      192 : rom_o = 12'b100100110100; //1.900000
      193 : rom_o = 12'b100100110100; //1.900000
      194 : rom_o = 12'b100100110100; //1.900000
      195 : rom_o = 12'b100100110100; //1.900000
      196 : rom_o = 12'b100100110100; //1.900000
      197 : rom_o = 12'b100100110100; //1.900000
      198 : rom_o = 12'b100100110100; //1.900000
      199 : rom_o = 12'b100100110100; //1.900000
      200 : rom_o = 12'b100110110000; //2.000000
      201 : rom_o = 12'b100110110000; //2.000000
      202 : rom_o = 12'b100110110000; //2.000000
      203 : rom_o = 12'b100110110000; //2.000000
      204 : rom_o = 12'b100110110000; //2.000000
      205 : rom_o = 12'b100110110000; //2.000000
      206 : rom_o = 12'b100110110000; //2.000000
      207 : rom_o = 12'b100110110000; //2.000000
      208 : rom_o = 12'b100110110000; //2.000000
      209 : rom_o = 12'b100110110000; //2.000000
      210 : rom_o = 12'b101000101100; //2.100000
      211 : rom_o = 12'b101000101100; //2.100000
      212 : rom_o = 12'b101000101100; //2.100000
      213 : rom_o = 12'b101000101100; //2.100000
      214 : rom_o = 12'b101000101100; //2.100000
      215 : rom_o = 12'b101000101100; //2.100000
      216 : rom_o = 12'b101000101100; //2.100000
      217 : rom_o = 12'b101000101100; //2.100000
      218 : rom_o = 12'b101000101100; //2.100000
      219 : rom_o = 12'b101000101100; //2.100000
      220 : rom_o = 12'b101010101000; //2.200000
      221 : rom_o = 12'b101010101000; //2.200000
      222 : rom_o = 12'b101010101000; //2.200000
      223 : rom_o = 12'b101010101000; //2.200000
      224 : rom_o = 12'b101010101000; //2.200000
      225 : rom_o = 12'b101010101000; //2.200000
      226 : rom_o = 12'b101010101000; //2.200000
      227 : rom_o = 12'b101010101000; //2.200000
      228 : rom_o = 12'b101010101000; //2.200000
      229 : rom_o = 12'b101010101000; //2.200000
      230 : rom_o = 12'b101100100100; //2.300000
      231 : rom_o = 12'b101100100100; //2.300000
      232 : rom_o = 12'b101100100100; //2.300000
      233 : rom_o = 12'b101100100100; //2.300000
      234 : rom_o = 12'b101100100100; //2.300000
      235 : rom_o = 12'b101100100100; //2.300000
      236 : rom_o = 12'b101100100100; //2.300000
      237 : rom_o = 12'b101100100100; //2.300000
      238 : rom_o = 12'b101100100100; //2.300000
      239 : rom_o = 12'b101100100100; //2.300000
      240 : rom_o = 12'b101110100000; //2.400000
      241 : rom_o = 12'b101110100000; //2.400000
      242 : rom_o = 12'b101110100000; //2.400000
      243 : rom_o = 12'b101110100000; //2.400000
      244 : rom_o = 12'b101110100000; //2.400000
      245 : rom_o = 12'b101110100000; //2.400000
      246 : rom_o = 12'b101110100000; //2.400000
      247 : rom_o = 12'b101110100000; //2.400000
      248 : rom_o = 12'b101110100000; //2.400000
      249 : rom_o = 12'b101110100000; //2.400000
      250 : rom_o = 12'b110000011100; //2.500000
      251 : rom_o = 12'b110000011100; //2.500000
      252 : rom_o = 12'b110000011100; //2.500000
      253 : rom_o = 12'b110000011100; //2.500000
      254 : rom_o = 12'b110000011100; //2.500000
      255 : rom_o = 12'b110000011100; //2.500000
      256 : rom_o = 12'b110000011100; //2.500000
      257 : rom_o = 12'b110000011100; //2.500000
      258 : rom_o = 12'b110000011100; //2.500000
      259 : rom_o = 12'b110000011100; //2.500000
      260 : rom_o = 12'b110010011000; //2.600000
      261 : rom_o = 12'b110010011000; //2.600000
      262 : rom_o = 12'b110010011000; //2.600000
      263 : rom_o = 12'b110010011000; //2.600000
      264 : rom_o = 12'b110010011000; //2.600000
      265 : rom_o = 12'b110010011000; //2.600000
      266 : rom_o = 12'b110010011000; //2.600000
      267 : rom_o = 12'b110010011000; //2.600000
      268 : rom_o = 12'b110010011000; //2.600000
      269 : rom_o = 12'b110010011000; //2.600000
      270 : rom_o = 12'b110100010100; //2.700000
      271 : rom_o = 12'b110100010100; //2.700000
      272 : rom_o = 12'b110100010100; //2.700000
      273 : rom_o = 12'b110100010100; //2.700000
      274 : rom_o = 12'b110100010100; //2.700000
      275 : rom_o = 12'b110100010100; //2.700000
      276 : rom_o = 12'b110100010100; //2.700000
      277 : rom_o = 12'b110100010100; //2.700000
      278 : rom_o = 12'b110100010100; //2.700000
      279 : rom_o = 12'b110100010100; //2.700000
      280 : rom_o = 12'b110110010000; //2.800000
      281 : rom_o = 12'b110110010000; //2.800000
      282 : rom_o = 12'b110110010000; //2.800000
      283 : rom_o = 12'b110110010000; //2.800000
      284 : rom_o = 12'b110110010000; //2.800000
      285 : rom_o = 12'b110110010000; //2.800000
      286 : rom_o = 12'b110110010000; //2.800000
      287 : rom_o = 12'b110110010000; //2.800000
      288 : rom_o = 12'b110110010000; //2.800000
      289 : rom_o = 12'b110110010000; //2.800000
      290 : rom_o = 12'b111000001100; //2.900000
      291 : rom_o = 12'b111000001100; //2.900000
      292 : rom_o = 12'b111000001100; //2.900000
      293 : rom_o = 12'b111000001100; //2.900000
      294 : rom_o = 12'b111000001100; //2.900000
      295 : rom_o = 12'b111000001100; //2.900000
      296 : rom_o = 12'b111000001100; //2.900000
      297 : rom_o = 12'b111000001100; //2.900000
      298 : rom_o = 12'b111000001100; //2.900000
      299 : rom_o = 12'b111000001100; //2.900000
      300 : rom_o = 12'b111010001000; //3.000000
      301 : rom_o = 12'b111010001000; //3.000000
      302 : rom_o = 12'b111010001000; //3.000000
      303 : rom_o = 12'b111010001000; //3.000000
      304 : rom_o = 12'b111010001000; //3.000000
      305 : rom_o = 12'b111010001000; //3.000000
      306 : rom_o = 12'b111010001000; //3.000000
      307 : rom_o = 12'b111010001000; //3.000000
      308 : rom_o = 12'b111010001000; //3.000000
      309 : rom_o = 12'b111010001000; //3.000000  
	  default: rom_o = 12'b000000000000;
	endcase
endmodule