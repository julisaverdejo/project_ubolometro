// Author: Julisa Verdejo Palacios
// Name: rom_volts.v
//
// Description: 


module rom_volts (
  input      [9:0] addr_i,
  output reg [11:0] rom_o
);

  always@(addr_i)  
    case(addr_i)
        0 : rom_o = 12'b000000000000; //0.000000
        1 : rom_o = 12'b000000000000; //0.000000
        2 : rom_o = 12'b000000000000; //0.000000
        3 : rom_o = 12'b000000000000; //0.000000
        4 : rom_o = 12'b000000000000; //0.000000
        5 : rom_o = 12'b000000000000; //0.000000
        6 : rom_o = 12'b000000000000; //0.000000
        7 : rom_o = 12'b000000000000; //0.000000
        8 : rom_o = 12'b000000000000; //0.000000
        9 : rom_o = 12'b000000000000; //0.000000
       10 : rom_o = 12'b000000101101; //0.036264
       11 : rom_o = 12'b000000101101; //0.036264
       12 : rom_o = 12'b000000101101; //0.036264
       13 : rom_o = 12'b000000101101; //0.036264
       14 : rom_o = 12'b000000101101; //0.036264
       15 : rom_o = 12'b000000101101; //0.036264
       16 : rom_o = 12'b000000101101; //0.036264
       17 : rom_o = 12'b000000101101; //0.036264
       18 : rom_o = 12'b000000101101; //0.036264
       19 : rom_o = 12'b000000101101; //0.036264
       20 : rom_o = 12'b000001011010; //0.072527
       21 : rom_o = 12'b000001011010; //0.072527
       22 : rom_o = 12'b000001011010; //0.072527
       23 : rom_o = 12'b000001011010; //0.072527
       24 : rom_o = 12'b000001011010; //0.072527
       25 : rom_o = 12'b000001011010; //0.072527
       26 : rom_o = 12'b000001011010; //0.072527
       27 : rom_o = 12'b000001011010; //0.072527
       28 : rom_o = 12'b000001011010; //0.072527
       29 : rom_o = 12'b000001011010; //0.072527
       30 : rom_o = 12'b000010000111; //0.108791
       31 : rom_o = 12'b000010000111; //0.108791
       32 : rom_o = 12'b000010000111; //0.108791
       33 : rom_o = 12'b000010000111; //0.108791
       34 : rom_o = 12'b000010000111; //0.108791
       35 : rom_o = 12'b000010000111; //0.108791
       36 : rom_o = 12'b000010000111; //0.108791
       37 : rom_o = 12'b000010000111; //0.108791
       38 : rom_o = 12'b000010000111; //0.108791
       39 : rom_o = 12'b000010000111; //0.108791
       40 : rom_o = 12'b000010110100; //0.145055
       41 : rom_o = 12'b000010110100; //0.145055
       42 : rom_o = 12'b000010110100; //0.145055
       43 : rom_o = 12'b000010110100; //0.145055
       44 : rom_o = 12'b000010110100; //0.145055
       45 : rom_o = 12'b000010110100; //0.145055
       46 : rom_o = 12'b000010110100; //0.145055
       47 : rom_o = 12'b000010110100; //0.145055
       48 : rom_o = 12'b000010110100; //0.145055
       49 : rom_o = 12'b000010110100; //0.145055
       50 : rom_o = 12'b000011100001; //0.181319
       51 : rom_o = 12'b000011100001; //0.181319
       52 : rom_o = 12'b000011100001; //0.181319
       53 : rom_o = 12'b000011100001; //0.181319
       54 : rom_o = 12'b000011100001; //0.181319
       55 : rom_o = 12'b000011100001; //0.181319
       56 : rom_o = 12'b000011100001; //0.181319
       57 : rom_o = 12'b000011100001; //0.181319
       58 : rom_o = 12'b000011100001; //0.181319
       59 : rom_o = 12'b000011100001; //0.181319
       60 : rom_o = 12'b000100001110; //0.217582
       61 : rom_o = 12'b000100001110; //0.217582
       62 : rom_o = 12'b000100001110; //0.217582
       63 : rom_o = 12'b000100001110; //0.217582
       64 : rom_o = 12'b000100001110; //0.217582
       65 : rom_o = 12'b000100001110; //0.217582
       66 : rom_o = 12'b000100001110; //0.217582
       67 : rom_o = 12'b000100001110; //0.217582
       68 : rom_o = 12'b000100001110; //0.217582
       69 : rom_o = 12'b000100001110; //0.217582
       70 : rom_o = 12'b000100111011; //0.253846
       71 : rom_o = 12'b000100111011; //0.253846
       72 : rom_o = 12'b000100111011; //0.253846
       73 : rom_o = 12'b000100111011; //0.253846
       74 : rom_o = 12'b000100111011; //0.253846
       75 : rom_o = 12'b000100111011; //0.253846
       76 : rom_o = 12'b000100111011; //0.253846
       77 : rom_o = 12'b000100111011; //0.253846
       78 : rom_o = 12'b000100111011; //0.253846
       79 : rom_o = 12'b000100111011; //0.253846
       80 : rom_o = 12'b000101101000; //0.290110
       81 : rom_o = 12'b000101101000; //0.290110
       82 : rom_o = 12'b000101101000; //0.290110
       83 : rom_o = 12'b000101101000; //0.290110
       84 : rom_o = 12'b000101101000; //0.290110
       85 : rom_o = 12'b000101101000; //0.290110
       86 : rom_o = 12'b000101101000; //0.290110
       87 : rom_o = 12'b000101101000; //0.290110
       88 : rom_o = 12'b000101101000; //0.290110
       89 : rom_o = 12'b000101101000; //0.290110
       90 : rom_o = 12'b000110010101; //0.326374
       91 : rom_o = 12'b000110010101; //0.326374
       92 : rom_o = 12'b000110010101; //0.326374
       93 : rom_o = 12'b000110010101; //0.326374
       94 : rom_o = 12'b000110010101; //0.326374
       95 : rom_o = 12'b000110010101; //0.326374
       96 : rom_o = 12'b000110010101; //0.326374
       97 : rom_o = 12'b000110010101; //0.326374
       98 : rom_o = 12'b000110010101; //0.326374
       99 : rom_o = 12'b000110010101; //0.326374
      100 : rom_o = 12'b000111000010; //0.362637
      101 : rom_o = 12'b000111000010; //0.362637
      102 : rom_o = 12'b000111000010; //0.362637
      103 : rom_o = 12'b000111000010; //0.362637
      104 : rom_o = 12'b000111000010; //0.362637
      105 : rom_o = 12'b000111000010; //0.362637
      106 : rom_o = 12'b000111000010; //0.362637
      107 : rom_o = 12'b000111000010; //0.362637
      108 : rom_o = 12'b000111000010; //0.362637
      109 : rom_o = 12'b000111000010; //0.362637
      110 : rom_o = 12'b000111101111; //0.398901
      111 : rom_o = 12'b000111101111; //0.398901
      112 : rom_o = 12'b000111101111; //0.398901
      113 : rom_o = 12'b000111101111; //0.398901
      114 : rom_o = 12'b000111101111; //0.398901
      115 : rom_o = 12'b000111101111; //0.398901
      116 : rom_o = 12'b000111101111; //0.398901
      117 : rom_o = 12'b000111101111; //0.398901
      118 : rom_o = 12'b000111101111; //0.398901
      119 : rom_o = 12'b000111101111; //0.398901
      120 : rom_o = 12'b001000011100; //0.435165
      121 : rom_o = 12'b001000011100; //0.435165
      122 : rom_o = 12'b001000011100; //0.435165
      123 : rom_o = 12'b001000011100; //0.435165
      124 : rom_o = 12'b001000011100; //0.435165
      125 : rom_o = 12'b001000011100; //0.435165
      126 : rom_o = 12'b001000011100; //0.435165
      127 : rom_o = 12'b001000011100; //0.435165
      128 : rom_o = 12'b001000011100; //0.435165
      129 : rom_o = 12'b001000011100; //0.435165
      130 : rom_o = 12'b001001001001; //0.471429
      131 : rom_o = 12'b001001001001; //0.471429
      132 : rom_o = 12'b001001001001; //0.471429
      133 : rom_o = 12'b001001001001; //0.471429
      134 : rom_o = 12'b001001001001; //0.471429
      135 : rom_o = 12'b001001001001; //0.471429
      136 : rom_o = 12'b001001001001; //0.471429
      137 : rom_o = 12'b001001001001; //0.471429
      138 : rom_o = 12'b001001001001; //0.471429
      139 : rom_o = 12'b001001001001; //0.471429
      140 : rom_o = 12'b001001110110; //0.507692
      141 : rom_o = 12'b001001110110; //0.507692
      142 : rom_o = 12'b001001110110; //0.507692
      143 : rom_o = 12'b001001110110; //0.507692
      144 : rom_o = 12'b001001110110; //0.507692
      145 : rom_o = 12'b001001110110; //0.507692
      146 : rom_o = 12'b001001110110; //0.507692
      147 : rom_o = 12'b001001110110; //0.507692
      148 : rom_o = 12'b001001110110; //0.507692
      149 : rom_o = 12'b001001110110; //0.507692
      150 : rom_o = 12'b001010100011; //0.543956
      151 : rom_o = 12'b001010100011; //0.543956
      152 : rom_o = 12'b001010100011; //0.543956
      153 : rom_o = 12'b001010100011; //0.543956
      154 : rom_o = 12'b001010100011; //0.543956
      155 : rom_o = 12'b001010100011; //0.543956
      156 : rom_o = 12'b001010100011; //0.543956
      157 : rom_o = 12'b001010100011; //0.543956
      158 : rom_o = 12'b001010100011; //0.543956
      159 : rom_o = 12'b001010100011; //0.543956
      160 : rom_o = 12'b001011010000; //0.580220
      161 : rom_o = 12'b001011010000; //0.580220
      162 : rom_o = 12'b001011010000; //0.580220
      163 : rom_o = 12'b001011010000; //0.580220
      164 : rom_o = 12'b001011010000; //0.580220
      165 : rom_o = 12'b001011010000; //0.580220
      166 : rom_o = 12'b001011010000; //0.580220
      167 : rom_o = 12'b001011010000; //0.580220
      168 : rom_o = 12'b001011010000; //0.580220
      169 : rom_o = 12'b001011010000; //0.580220
      170 : rom_o = 12'b001011111101; //0.616484
      171 : rom_o = 12'b001011111101; //0.616484
      172 : rom_o = 12'b001011111101; //0.616484
      173 : rom_o = 12'b001011111101; //0.616484
      174 : rom_o = 12'b001011111101; //0.616484
      175 : rom_o = 12'b001011111101; //0.616484
      176 : rom_o = 12'b001011111101; //0.616484
      177 : rom_o = 12'b001011111101; //0.616484
      178 : rom_o = 12'b001011111101; //0.616484
      179 : rom_o = 12'b001011111101; //0.616484
      180 : rom_o = 12'b001100101010; //0.652747
      181 : rom_o = 12'b001100101010; //0.652747
      182 : rom_o = 12'b001100101010; //0.652747
      183 : rom_o = 12'b001100101010; //0.652747
      184 : rom_o = 12'b001100101010; //0.652747
      185 : rom_o = 12'b001100101010; //0.652747
      186 : rom_o = 12'b001100101010; //0.652747
      187 : rom_o = 12'b001100101010; //0.652747
      188 : rom_o = 12'b001100101010; //0.652747
      189 : rom_o = 12'b001100101010; //0.652747
      190 : rom_o = 12'b001101010111; //0.689011
      191 : rom_o = 12'b001101010111; //0.689011
      192 : rom_o = 12'b001101010111; //0.689011
      193 : rom_o = 12'b001101010111; //0.689011
      194 : rom_o = 12'b001101010111; //0.689011
      195 : rom_o = 12'b001101010111; //0.689011
      196 : rom_o = 12'b001101010111; //0.689011
      197 : rom_o = 12'b001101010111; //0.689011
      198 : rom_o = 12'b001101010111; //0.689011
      199 : rom_o = 12'b001101010111; //0.689011
      200 : rom_o = 12'b001110000100; //0.725275
      201 : rom_o = 12'b001110000100; //0.725275
      202 : rom_o = 12'b001110000100; //0.725275
      203 : rom_o = 12'b001110000100; //0.725275
      204 : rom_o = 12'b001110000100; //0.725275
      205 : rom_o = 12'b001110000100; //0.725275
      206 : rom_o = 12'b001110000100; //0.725275
      207 : rom_o = 12'b001110000100; //0.725275
      208 : rom_o = 12'b001110000100; //0.725275
      209 : rom_o = 12'b001110000100; //0.725275
      210 : rom_o = 12'b001110110001; //0.761538
      211 : rom_o = 12'b001110110001; //0.761538
      212 : rom_o = 12'b001110110001; //0.761538
      213 : rom_o = 12'b001110110001; //0.761538
      214 : rom_o = 12'b001110110001; //0.761538
      215 : rom_o = 12'b001110110001; //0.761538
      216 : rom_o = 12'b001110110001; //0.761538
      217 : rom_o = 12'b001110110001; //0.761538
      218 : rom_o = 12'b001110110001; //0.761538
      219 : rom_o = 12'b001110110001; //0.761538
      220 : rom_o = 12'b001111011110; //0.797802
      221 : rom_o = 12'b001111011110; //0.797802
      222 : rom_o = 12'b001111011110; //0.797802
      223 : rom_o = 12'b001111011110; //0.797802
      224 : rom_o = 12'b001111011110; //0.797802
      225 : rom_o = 12'b001111011110; //0.797802
      226 : rom_o = 12'b001111011110; //0.797802
      227 : rom_o = 12'b001111011110; //0.797802
      228 : rom_o = 12'b001111011110; //0.797802
      229 : rom_o = 12'b001111011110; //0.797802
      230 : rom_o = 12'b010000001011; //0.834066
      231 : rom_o = 12'b010000001011; //0.834066
      232 : rom_o = 12'b010000001011; //0.834066
      233 : rom_o = 12'b010000001011; //0.834066
      234 : rom_o = 12'b010000001011; //0.834066
      235 : rom_o = 12'b010000001011; //0.834066
      236 : rom_o = 12'b010000001011; //0.834066
      237 : rom_o = 12'b010000001011; //0.834066
      238 : rom_o = 12'b010000001011; //0.834066
      239 : rom_o = 12'b010000001011; //0.834066
      240 : rom_o = 12'b010000111000; //0.870330
      241 : rom_o = 12'b010000111000; //0.870330
      242 : rom_o = 12'b010000111000; //0.870330
      243 : rom_o = 12'b010000111000; //0.870330
      244 : rom_o = 12'b010000111000; //0.870330
      245 : rom_o = 12'b010000111000; //0.870330
      246 : rom_o = 12'b010000111000; //0.870330
      247 : rom_o = 12'b010000111000; //0.870330
      248 : rom_o = 12'b010000111000; //0.870330
      249 : rom_o = 12'b010000111000; //0.870330
      250 : rom_o = 12'b010001100101; //0.906593
      251 : rom_o = 12'b010001100101; //0.906593
      252 : rom_o = 12'b010001100101; //0.906593
      253 : rom_o = 12'b010001100101; //0.906593
      254 : rom_o = 12'b010001100101; //0.906593
      255 : rom_o = 12'b010001100101; //0.906593
      256 : rom_o = 12'b010001100101; //0.906593
      257 : rom_o = 12'b010001100101; //0.906593
      258 : rom_o = 12'b010001100101; //0.906593
      259 : rom_o = 12'b010001100101; //0.906593
      260 : rom_o = 12'b010010010010; //0.942857
      261 : rom_o = 12'b010010010010; //0.942857
      262 : rom_o = 12'b010010010010; //0.942857
      263 : rom_o = 12'b010010010010; //0.942857
      264 : rom_o = 12'b010010010010; //0.942857
      265 : rom_o = 12'b010010010010; //0.942857
      266 : rom_o = 12'b010010010010; //0.942857
      267 : rom_o = 12'b010010010010; //0.942857
      268 : rom_o = 12'b010010010010; //0.942857
      269 : rom_o = 12'b010010010010; //0.942857
      270 : rom_o = 12'b010010111111; //0.979121
      271 : rom_o = 12'b010010111111; //0.979121
      272 : rom_o = 12'b010010111111; //0.979121
      273 : rom_o = 12'b010010111111; //0.979121
      274 : rom_o = 12'b010010111111; //0.979121
      275 : rom_o = 12'b010010111111; //0.979121
      276 : rom_o = 12'b010010111111; //0.979121
      277 : rom_o = 12'b010010111111; //0.979121
      278 : rom_o = 12'b010010111111; //0.979121
      279 : rom_o = 12'b010010111111; //0.979121
      280 : rom_o = 12'b010011101100; //1.015385
      281 : rom_o = 12'b010011101100; //1.015385
      282 : rom_o = 12'b010011101100; //1.015385
      283 : rom_o = 12'b010011101100; //1.015385
      284 : rom_o = 12'b010011101100; //1.015385
      285 : rom_o = 12'b010011101100; //1.015385
      286 : rom_o = 12'b010011101100; //1.015385
      287 : rom_o = 12'b010011101100; //1.015385
      288 : rom_o = 12'b010011101100; //1.015385
      289 : rom_o = 12'b010011101100; //1.015385
      290 : rom_o = 12'b010100011001; //1.051648
      291 : rom_o = 12'b010100011001; //1.051648
      292 : rom_o = 12'b010100011001; //1.051648
      293 : rom_o = 12'b010100011001; //1.051648
      294 : rom_o = 12'b010100011001; //1.051648
      295 : rom_o = 12'b010100011001; //1.051648
      296 : rom_o = 12'b010100011001; //1.051648
      297 : rom_o = 12'b010100011001; //1.051648
      298 : rom_o = 12'b010100011001; //1.051648
      299 : rom_o = 12'b010100011001; //1.051648
      300 : rom_o = 12'b010101000110; //1.087912
      301 : rom_o = 12'b010101000110; //1.087912
      302 : rom_o = 12'b010101000110; //1.087912
      303 : rom_o = 12'b010101000110; //1.087912
      304 : rom_o = 12'b010101000110; //1.087912
      305 : rom_o = 12'b010101000110; //1.087912
      306 : rom_o = 12'b010101000110; //1.087912
      307 : rom_o = 12'b010101000110; //1.087912
      308 : rom_o = 12'b010101000110; //1.087912
      309 : rom_o = 12'b010101000110; //1.087912
      310 : rom_o = 12'b010101110011; //1.124176
      311 : rom_o = 12'b010101110011; //1.124176
      312 : rom_o = 12'b010101110011; //1.124176
      313 : rom_o = 12'b010101110011; //1.124176
      314 : rom_o = 12'b010101110011; //1.124176
      315 : rom_o = 12'b010101110011; //1.124176
      316 : rom_o = 12'b010101110011; //1.124176
      317 : rom_o = 12'b010101110011; //1.124176
      318 : rom_o = 12'b010101110011; //1.124176
      319 : rom_o = 12'b010101110011; //1.124176
      320 : rom_o = 12'b010110100000; //1.160440
      321 : rom_o = 12'b010110100000; //1.160440
      322 : rom_o = 12'b010110100000; //1.160440
      323 : rom_o = 12'b010110100000; //1.160440
      324 : rom_o = 12'b010110100000; //1.160440
      325 : rom_o = 12'b010110100000; //1.160440
      326 : rom_o = 12'b010110100000; //1.160440
      327 : rom_o = 12'b010110100000; //1.160440
      328 : rom_o = 12'b010110100000; //1.160440
      329 : rom_o = 12'b010110100000; //1.160440
      330 : rom_o = 12'b010111001101; //1.196703
      331 : rom_o = 12'b010111001101; //1.196703
      332 : rom_o = 12'b010111001101; //1.196703
      333 : rom_o = 12'b010111001101; //1.196703
      334 : rom_o = 12'b010111001101; //1.196703
      335 : rom_o = 12'b010111001101; //1.196703
      336 : rom_o = 12'b010111001101; //1.196703
      337 : rom_o = 12'b010111001101; //1.196703
      338 : rom_o = 12'b010111001101; //1.196703
      339 : rom_o = 12'b010111001101; //1.196703
      340 : rom_o = 12'b010111111010; //1.232967
      341 : rom_o = 12'b010111111010; //1.232967
      342 : rom_o = 12'b010111111010; //1.232967
      343 : rom_o = 12'b010111111010; //1.232967
      344 : rom_o = 12'b010111111010; //1.232967
      345 : rom_o = 12'b010111111010; //1.232967
      346 : rom_o = 12'b010111111010; //1.232967
      347 : rom_o = 12'b010111111010; //1.232967
      348 : rom_o = 12'b010111111010; //1.232967
      349 : rom_o = 12'b010111111010; //1.232967
      350 : rom_o = 12'b011000100111; //1.269231
      351 : rom_o = 12'b011000100111; //1.269231
      352 : rom_o = 12'b011000100111; //1.269231
      353 : rom_o = 12'b011000100111; //1.269231
      354 : rom_o = 12'b011000100111; //1.269231
      355 : rom_o = 12'b011000100111; //1.269231
      356 : rom_o = 12'b011000100111; //1.269231
      357 : rom_o = 12'b011000100111; //1.269231
      358 : rom_o = 12'b011000100111; //1.269231
      359 : rom_o = 12'b011000100111; //1.269231
      360 : rom_o = 12'b011001010100; //1.305495
      361 : rom_o = 12'b011001010100; //1.305495
      362 : rom_o = 12'b011001010100; //1.305495
      363 : rom_o = 12'b011001010100; //1.305495
      364 : rom_o = 12'b011001010100; //1.305495
      365 : rom_o = 12'b011001010100; //1.305495
      366 : rom_o = 12'b011001010100; //1.305495
      367 : rom_o = 12'b011001010100; //1.305495
      368 : rom_o = 12'b011001010100; //1.305495
      369 : rom_o = 12'b011001010100; //1.305495
      370 : rom_o = 12'b011010000001; //1.341758
      371 : rom_o = 12'b011010000001; //1.341758
      372 : rom_o = 12'b011010000001; //1.341758
      373 : rom_o = 12'b011010000001; //1.341758
      374 : rom_o = 12'b011010000001; //1.341758
      375 : rom_o = 12'b011010000001; //1.341758
      376 : rom_o = 12'b011010000001; //1.341758
      377 : rom_o = 12'b011010000001; //1.341758
      378 : rom_o = 12'b011010000001; //1.341758
      379 : rom_o = 12'b011010000001; //1.341758
      380 : rom_o = 12'b011010101110; //1.378022
      381 : rom_o = 12'b011010101110; //1.378022
      382 : rom_o = 12'b011010101110; //1.378022
      383 : rom_o = 12'b011010101110; //1.378022
      384 : rom_o = 12'b011010101110; //1.378022
      385 : rom_o = 12'b011010101110; //1.378022
      386 : rom_o = 12'b011010101110; //1.378022
      387 : rom_o = 12'b011010101110; //1.378022
      388 : rom_o = 12'b011010101110; //1.378022
      389 : rom_o = 12'b011010101110; //1.378022
      390 : rom_o = 12'b011011011011; //1.414286
      391 : rom_o = 12'b011011011011; //1.414286
      392 : rom_o = 12'b011011011011; //1.414286
      393 : rom_o = 12'b011011011011; //1.414286
      394 : rom_o = 12'b011011011011; //1.414286
      395 : rom_o = 12'b011011011011; //1.414286
      396 : rom_o = 12'b011011011011; //1.414286
      397 : rom_o = 12'b011011011011; //1.414286
      398 : rom_o = 12'b011011011011; //1.414286
      399 : rom_o = 12'b011011011011; //1.414286
      400 : rom_o = 12'b011100001000; //1.450549
      401 : rom_o = 12'b011100001000; //1.450549
      402 : rom_o = 12'b011100001000; //1.450549
      403 : rom_o = 12'b011100001000; //1.450549
      404 : rom_o = 12'b011100001000; //1.450549
      405 : rom_o = 12'b011100001000; //1.450549
      406 : rom_o = 12'b011100001000; //1.450549
      407 : rom_o = 12'b011100001000; //1.450549
      408 : rom_o = 12'b011100001000; //1.450549
      409 : rom_o = 12'b011100001000; //1.450549
      410 : rom_o = 12'b011100110101; //1.486813
      411 : rom_o = 12'b011100110101; //1.486813
      412 : rom_o = 12'b011100110101; //1.486813
      413 : rom_o = 12'b011100110101; //1.486813
      414 : rom_o = 12'b011100110101; //1.486813
      415 : rom_o = 12'b011100110101; //1.486813
      416 : rom_o = 12'b011100110101; //1.486813
      417 : rom_o = 12'b011100110101; //1.486813
      418 : rom_o = 12'b011100110101; //1.486813
      419 : rom_o = 12'b011100110101; //1.486813
      420 : rom_o = 12'b011101100010; //1.523077
      421 : rom_o = 12'b011101100010; //1.523077
      422 : rom_o = 12'b011101100010; //1.523077
      423 : rom_o = 12'b011101100010; //1.523077
      424 : rom_o = 12'b011101100010; //1.523077
      425 : rom_o = 12'b011101100010; //1.523077
      426 : rom_o = 12'b011101100010; //1.523077
      427 : rom_o = 12'b011101100010; //1.523077
      428 : rom_o = 12'b011101100010; //1.523077
      429 : rom_o = 12'b011101100010; //1.523077
      430 : rom_o = 12'b011110001111; //1.559341
      431 : rom_o = 12'b011110001111; //1.559341
      432 : rom_o = 12'b011110001111; //1.559341
      433 : rom_o = 12'b011110001111; //1.559341
      434 : rom_o = 12'b011110001111; //1.559341
      435 : rom_o = 12'b011110001111; //1.559341
      436 : rom_o = 12'b011110001111; //1.559341
      437 : rom_o = 12'b011110001111; //1.559341
      438 : rom_o = 12'b011110001111; //1.559341
      439 : rom_o = 12'b011110001111; //1.559341
      440 : rom_o = 12'b011110111100; //1.595604
      441 : rom_o = 12'b011110111100; //1.595604
      442 : rom_o = 12'b011110111100; //1.595604
      443 : rom_o = 12'b011110111100; //1.595604
      444 : rom_o = 12'b011110111100; //1.595604
      445 : rom_o = 12'b011110111100; //1.595604
      446 : rom_o = 12'b011110111100; //1.595604
      447 : rom_o = 12'b011110111100; //1.595604
      448 : rom_o = 12'b011110111100; //1.595604
      449 : rom_o = 12'b011110111100; //1.595604
      450 : rom_o = 12'b011111101001; //1.631868
      451 : rom_o = 12'b011111101001; //1.631868
      452 : rom_o = 12'b011111101001; //1.631868
      453 : rom_o = 12'b011111101001; //1.631868
      454 : rom_o = 12'b011111101001; //1.631868
      455 : rom_o = 12'b011111101001; //1.631868
      456 : rom_o = 12'b011111101001; //1.631868
      457 : rom_o = 12'b011111101001; //1.631868
      458 : rom_o = 12'b011111101001; //1.631868
      459 : rom_o = 12'b011111101001; //1.631868
      460 : rom_o = 12'b100000010110; //1.668132
      461 : rom_o = 12'b100000010110; //1.668132
      462 : rom_o = 12'b100000010110; //1.668132
      463 : rom_o = 12'b100000010110; //1.668132
      464 : rom_o = 12'b100000010110; //1.668132
      465 : rom_o = 12'b100000010110; //1.668132
      466 : rom_o = 12'b100000010110; //1.668132
      467 : rom_o = 12'b100000010110; //1.668132
      468 : rom_o = 12'b100000010110; //1.668132
      469 : rom_o = 12'b100000010110; //1.668132
      470 : rom_o = 12'b100001000011; //1.704396
      471 : rom_o = 12'b100001000011; //1.704396
      472 : rom_o = 12'b100001000011; //1.704396
      473 : rom_o = 12'b100001000011; //1.704396
      474 : rom_o = 12'b100001000011; //1.704396
      475 : rom_o = 12'b100001000011; //1.704396
      476 : rom_o = 12'b100001000011; //1.704396
      477 : rom_o = 12'b100001000011; //1.704396
      478 : rom_o = 12'b100001000011; //1.704396
      479 : rom_o = 12'b100001000011; //1.704396
      480 : rom_o = 12'b100001110000; //1.740659
      481 : rom_o = 12'b100001110000; //1.740659
      482 : rom_o = 12'b100001110000; //1.740659
      483 : rom_o = 12'b100001110000; //1.740659
      484 : rom_o = 12'b100001110000; //1.740659
      485 : rom_o = 12'b100001110000; //1.740659
      486 : rom_o = 12'b100001110000; //1.740659
      487 : rom_o = 12'b100001110000; //1.740659
      488 : rom_o = 12'b100001110000; //1.740659
      489 : rom_o = 12'b100001110000; //1.740659
      490 : rom_o = 12'b100010011101; //1.776923
      491 : rom_o = 12'b100010011101; //1.776923
      492 : rom_o = 12'b100010011101; //1.776923
      493 : rom_o = 12'b100010011101; //1.776923
      494 : rom_o = 12'b100010011101; //1.776923
      495 : rom_o = 12'b100010011101; //1.776923
      496 : rom_o = 12'b100010011101; //1.776923
      497 : rom_o = 12'b100010011101; //1.776923
      498 : rom_o = 12'b100010011101; //1.776923
      499 : rom_o = 12'b100010011101; //1.776923
      500 : rom_o = 12'b100011001010; //1.813187
      501 : rom_o = 12'b100011001010; //1.813187
      502 : rom_o = 12'b100011001010; //1.813187
      503 : rom_o = 12'b100011001010; //1.813187
      504 : rom_o = 12'b100011001010; //1.813187
      505 : rom_o = 12'b100011001010; //1.813187
      506 : rom_o = 12'b100011001010; //1.813187
      507 : rom_o = 12'b100011001010; //1.813187
      508 : rom_o = 12'b100011001010; //1.813187
      509 : rom_o = 12'b100011001010; //1.813187
      510 : rom_o = 12'b100011110111; //1.849451
      511 : rom_o = 12'b100011110111; //1.849451
      512 : rom_o = 12'b100011110111; //1.849451
      513 : rom_o = 12'b100011110111; //1.849451
      514 : rom_o = 12'b100011110111; //1.849451
      515 : rom_o = 12'b100011110111; //1.849451
      516 : rom_o = 12'b100011110111; //1.849451
      517 : rom_o = 12'b100011110111; //1.849451
      518 : rom_o = 12'b100011110111; //1.849451
      519 : rom_o = 12'b100011110111; //1.849451
      520 : rom_o = 12'b100100100100; //1.885714
      521 : rom_o = 12'b100100100100; //1.885714
      522 : rom_o = 12'b100100100100; //1.885714
      523 : rom_o = 12'b100100100100; //1.885714
      524 : rom_o = 12'b100100100100; //1.885714
      525 : rom_o = 12'b100100100100; //1.885714
      526 : rom_o = 12'b100100100100; //1.885714
      527 : rom_o = 12'b100100100100; //1.885714
      528 : rom_o = 12'b100100100100; //1.885714
      529 : rom_o = 12'b100100100100; //1.885714
      530 : rom_o = 12'b100101010001; //1.921978
      531 : rom_o = 12'b100101010001; //1.921978
      532 : rom_o = 12'b100101010001; //1.921978
      533 : rom_o = 12'b100101010001; //1.921978
      534 : rom_o = 12'b100101010001; //1.921978
      535 : rom_o = 12'b100101010001; //1.921978
      536 : rom_o = 12'b100101010001; //1.921978
      537 : rom_o = 12'b100101010001; //1.921978
      538 : rom_o = 12'b100101010001; //1.921978
      539 : rom_o = 12'b100101010001; //1.921978
      540 : rom_o = 12'b100101111110; //1.958242
      541 : rom_o = 12'b100101111110; //1.958242
      542 : rom_o = 12'b100101111110; //1.958242
      543 : rom_o = 12'b100101111110; //1.958242
      544 : rom_o = 12'b100101111110; //1.958242
      545 : rom_o = 12'b100101111110; //1.958242
      546 : rom_o = 12'b100101111110; //1.958242
      547 : rom_o = 12'b100101111110; //1.958242
      548 : rom_o = 12'b100101111110; //1.958242
      549 : rom_o = 12'b100101111110; //1.958242
      550 : rom_o = 12'b100110101011; //1.994505
      551 : rom_o = 12'b100110101011; //1.994505
      552 : rom_o = 12'b100110101011; //1.994505
      553 : rom_o = 12'b100110101011; //1.994505
      554 : rom_o = 12'b100110101011; //1.994505
      555 : rom_o = 12'b100110101011; //1.994505
      556 : rom_o = 12'b100110101011; //1.994505
      557 : rom_o = 12'b100110101011; //1.994505
      558 : rom_o = 12'b100110101011; //1.994505
      559 : rom_o = 12'b100110101011; //1.994505
      560 : rom_o = 12'b100111011000; //2.030769
      561 : rom_o = 12'b100111011000; //2.030769
      562 : rom_o = 12'b100111011000; //2.030769
      563 : rom_o = 12'b100111011000; //2.030769
      564 : rom_o = 12'b100111011000; //2.030769
      565 : rom_o = 12'b100111011000; //2.030769
      566 : rom_o = 12'b100111011000; //2.030769
      567 : rom_o = 12'b100111011000; //2.030769
      568 : rom_o = 12'b100111011000; //2.030769
      569 : rom_o = 12'b100111011000; //2.030769
      570 : rom_o = 12'b101000000101; //2.067033
      571 : rom_o = 12'b101000000101; //2.067033
      572 : rom_o = 12'b101000000101; //2.067033
      573 : rom_o = 12'b101000000101; //2.067033
      574 : rom_o = 12'b101000000101; //2.067033
      575 : rom_o = 12'b101000000101; //2.067033
      576 : rom_o = 12'b101000000101; //2.067033
      577 : rom_o = 12'b101000000101; //2.067033
      578 : rom_o = 12'b101000000101; //2.067033
      579 : rom_o = 12'b101000000101; //2.067033
      580 : rom_o = 12'b101000110010; //2.103297
      581 : rom_o = 12'b101000110010; //2.103297
      582 : rom_o = 12'b101000110010; //2.103297
      583 : rom_o = 12'b101000110010; //2.103297
      584 : rom_o = 12'b101000110010; //2.103297
      585 : rom_o = 12'b101000110010; //2.103297
      586 : rom_o = 12'b101000110010; //2.103297
      587 : rom_o = 12'b101000110010; //2.103297
      588 : rom_o = 12'b101000110010; //2.103297
      589 : rom_o = 12'b101000110010; //2.103297
      590 : rom_o = 12'b101001011111; //2.139560
      591 : rom_o = 12'b101001011111; //2.139560
      592 : rom_o = 12'b101001011111; //2.139560
      593 : rom_o = 12'b101001011111; //2.139560
      594 : rom_o = 12'b101001011111; //2.139560
      595 : rom_o = 12'b101001011111; //2.139560
      596 : rom_o = 12'b101001011111; //2.139560
      597 : rom_o = 12'b101001011111; //2.139560
      598 : rom_o = 12'b101001011111; //2.139560
      599 : rom_o = 12'b101001011111; //2.139560
      600 : rom_o = 12'b101010001100; //2.175824
      601 : rom_o = 12'b101010001100; //2.175824
      602 : rom_o = 12'b101010001100; //2.175824
      603 : rom_o = 12'b101010001100; //2.175824
      604 : rom_o = 12'b101010001100; //2.175824
      605 : rom_o = 12'b101010001100; //2.175824
      606 : rom_o = 12'b101010001100; //2.175824
      607 : rom_o = 12'b101010001100; //2.175824
      608 : rom_o = 12'b101010001100; //2.175824
      609 : rom_o = 12'b101010001100; //2.175824
      610 : rom_o = 12'b101010111001; //2.212088
      611 : rom_o = 12'b101010111001; //2.212088
      612 : rom_o = 12'b101010111001; //2.212088
      613 : rom_o = 12'b101010111001; //2.212088
      614 : rom_o = 12'b101010111001; //2.212088
      615 : rom_o = 12'b101010111001; //2.212088
      616 : rom_o = 12'b101010111001; //2.212088
      617 : rom_o = 12'b101010111001; //2.212088
      618 : rom_o = 12'b101010111001; //2.212088
      619 : rom_o = 12'b101010111001; //2.212088
      620 : rom_o = 12'b101011100110; //2.248352
      621 : rom_o = 12'b101011100110; //2.248352
      622 : rom_o = 12'b101011100110; //2.248352
      623 : rom_o = 12'b101011100110; //2.248352
      624 : rom_o = 12'b101011100110; //2.248352
      625 : rom_o = 12'b101011100110; //2.248352
      626 : rom_o = 12'b101011100110; //2.248352
      627 : rom_o = 12'b101011100110; //2.248352
      628 : rom_o = 12'b101011100110; //2.248352
      629 : rom_o = 12'b101011100110; //2.248352
      630 : rom_o = 12'b101100010011; //2.284615
      631 : rom_o = 12'b101100010011; //2.284615
      632 : rom_o = 12'b101100010011; //2.284615
      633 : rom_o = 12'b101100010011; //2.284615
      634 : rom_o = 12'b101100010011; //2.284615
      635 : rom_o = 12'b101100010011; //2.284615
      636 : rom_o = 12'b101100010011; //2.284615
      637 : rom_o = 12'b101100010011; //2.284615
      638 : rom_o = 12'b101100010011; //2.284615
      639 : rom_o = 12'b101100010011; //2.284615
      640 : rom_o = 12'b101101000000; //2.320879
      641 : rom_o = 12'b101101000000; //2.320879
      642 : rom_o = 12'b101101000000; //2.320879
      643 : rom_o = 12'b101101000000; //2.320879
      644 : rom_o = 12'b101101000000; //2.320879
      645 : rom_o = 12'b101101000000; //2.320879
      646 : rom_o = 12'b101101000000; //2.320879
      647 : rom_o = 12'b101101000000; //2.320879
      648 : rom_o = 12'b101101000000; //2.320879
      649 : rom_o = 12'b101101000000; //2.320879
      650 : rom_o = 12'b101101101101; //2.357143
      651 : rom_o = 12'b101101101101; //2.357143
      652 : rom_o = 12'b101101101101; //2.357143
      653 : rom_o = 12'b101101101101; //2.357143
      654 : rom_o = 12'b101101101101; //2.357143
      655 : rom_o = 12'b101101101101; //2.357143
      656 : rom_o = 12'b101101101101; //2.357143
      657 : rom_o = 12'b101101101101; //2.357143
      658 : rom_o = 12'b101101101101; //2.357143
      659 : rom_o = 12'b101101101101; //2.357143
      660 : rom_o = 12'b101110011010; //2.393407
      661 : rom_o = 12'b101110011010; //2.393407
      662 : rom_o = 12'b101110011010; //2.393407
      663 : rom_o = 12'b101110011010; //2.393407
      664 : rom_o = 12'b101110011010; //2.393407
      665 : rom_o = 12'b101110011010; //2.393407
      666 : rom_o = 12'b101110011010; //2.393407
      667 : rom_o = 12'b101110011010; //2.393407
      668 : rom_o = 12'b101110011010; //2.393407
      669 : rom_o = 12'b101110011010; //2.393407
      670 : rom_o = 12'b101111000111; //2.429670
      671 : rom_o = 12'b101111000111; //2.429670
      672 : rom_o = 12'b101111000111; //2.429670
      673 : rom_o = 12'b101111000111; //2.429670
      674 : rom_o = 12'b101111000111; //2.429670
      675 : rom_o = 12'b101111000111; //2.429670
      676 : rom_o = 12'b101111000111; //2.429670
      677 : rom_o = 12'b101111000111; //2.429670
      678 : rom_o = 12'b101111000111; //2.429670
      679 : rom_o = 12'b101111000111; //2.429670
      680 : rom_o = 12'b101111110100; //2.465934
      681 : rom_o = 12'b101111110100; //2.465934
      682 : rom_o = 12'b101111110100; //2.465934
      683 : rom_o = 12'b101111110100; //2.465934
      684 : rom_o = 12'b101111110100; //2.465934
      685 : rom_o = 12'b101111110100; //2.465934
      686 : rom_o = 12'b101111110100; //2.465934
      687 : rom_o = 12'b101111110100; //2.465934
      688 : rom_o = 12'b101111110100; //2.465934
      689 : rom_o = 12'b101111110100; //2.465934
      690 : rom_o = 12'b110000100001; //2.502198
      691 : rom_o = 12'b110000100001; //2.502198
      692 : rom_o = 12'b110000100001; //2.502198
      693 : rom_o = 12'b110000100001; //2.502198
      694 : rom_o = 12'b110000100001; //2.502198
      695 : rom_o = 12'b110000100001; //2.502198
      696 : rom_o = 12'b110000100001; //2.502198
      697 : rom_o = 12'b110000100001; //2.502198
      698 : rom_o = 12'b110000100001; //2.502198
      699 : rom_o = 12'b110000100001; //2.502198
      700 : rom_o = 12'b110001001110; //2.538462
      701 : rom_o = 12'b110001001110; //2.538462
      702 : rom_o = 12'b110001001110; //2.538462
      703 : rom_o = 12'b110001001110; //2.538462
      704 : rom_o = 12'b110001001110; //2.538462
      705 : rom_o = 12'b110001001110; //2.538462
      706 : rom_o = 12'b110001001110; //2.538462
      707 : rom_o = 12'b110001001110; //2.538462
      708 : rom_o = 12'b110001001110; //2.538462
      709 : rom_o = 12'b110001001110; //2.538462
      710 : rom_o = 12'b110001111011; //2.574725
      711 : rom_o = 12'b110001111011; //2.574725
      712 : rom_o = 12'b110001111011; //2.574725
      713 : rom_o = 12'b110001111011; //2.574725
      714 : rom_o = 12'b110001111011; //2.574725
      715 : rom_o = 12'b110001111011; //2.574725
      716 : rom_o = 12'b110001111011; //2.574725
      717 : rom_o = 12'b110001111011; //2.574725
      718 : rom_o = 12'b110001111011; //2.574725
      719 : rom_o = 12'b110001111011; //2.574725
      720 : rom_o = 12'b110010101000; //2.610989
      721 : rom_o = 12'b110010101000; //2.610989
      722 : rom_o = 12'b110010101000; //2.610989
      723 : rom_o = 12'b110010101000; //2.610989
      724 : rom_o = 12'b110010101000; //2.610989
      725 : rom_o = 12'b110010101000; //2.610989
      726 : rom_o = 12'b110010101000; //2.610989
      727 : rom_o = 12'b110010101000; //2.610989
      728 : rom_o = 12'b110010101000; //2.610989
      729 : rom_o = 12'b110010101000; //2.610989
      730 : rom_o = 12'b110011010101; //2.647253
      731 : rom_o = 12'b110011010101; //2.647253
      732 : rom_o = 12'b110011010101; //2.647253
      733 : rom_o = 12'b110011010101; //2.647253
      734 : rom_o = 12'b110011010101; //2.647253
      735 : rom_o = 12'b110011010101; //2.647253
      736 : rom_o = 12'b110011010101; //2.647253
      737 : rom_o = 12'b110011010101; //2.647253
      738 : rom_o = 12'b110011010101; //2.647253
      739 : rom_o = 12'b110011010101; //2.647253
      740 : rom_o = 12'b110100000010; //2.683516
      741 : rom_o = 12'b110100000010; //2.683516
      742 : rom_o = 12'b110100000010; //2.683516
      743 : rom_o = 12'b110100000010; //2.683516
      744 : rom_o = 12'b110100000010; //2.683516
      745 : rom_o = 12'b110100000010; //2.683516
      746 : rom_o = 12'b110100000010; //2.683516
      747 : rom_o = 12'b110100000010; //2.683516
      748 : rom_o = 12'b110100000010; //2.683516
      749 : rom_o = 12'b110100000010; //2.683516
      750 : rom_o = 12'b110100101111; //2.719780
      751 : rom_o = 12'b110100101111; //2.719780
      752 : rom_o = 12'b110100101111; //2.719780
      753 : rom_o = 12'b110100101111; //2.719780
      754 : rom_o = 12'b110100101111; //2.719780
      755 : rom_o = 12'b110100101111; //2.719780
      756 : rom_o = 12'b110100101111; //2.719780
      757 : rom_o = 12'b110100101111; //2.719780
      758 : rom_o = 12'b110100101111; //2.719780
      759 : rom_o = 12'b110100101111; //2.719780
      760 : rom_o = 12'b110101011100; //2.756044
      761 : rom_o = 12'b110101011100; //2.756044
      762 : rom_o = 12'b110101011100; //2.756044
      763 : rom_o = 12'b110101011100; //2.756044
      764 : rom_o = 12'b110101011100; //2.756044
      765 : rom_o = 12'b110101011100; //2.756044
      766 : rom_o = 12'b110101011100; //2.756044
      767 : rom_o = 12'b110101011100; //2.756044
      768 : rom_o = 12'b110101011100; //2.756044
      769 : rom_o = 12'b110101011100; //2.756044
      770 : rom_o = 12'b110110001001; //2.792308
      771 : rom_o = 12'b110110001001; //2.792308
      772 : rom_o = 12'b110110001001; //2.792308
      773 : rom_o = 12'b110110001001; //2.792308
      774 : rom_o = 12'b110110001001; //2.792308
      775 : rom_o = 12'b110110001001; //2.792308
      776 : rom_o = 12'b110110001001; //2.792308
      777 : rom_o = 12'b110110001001; //2.792308
      778 : rom_o = 12'b110110001001; //2.792308
      779 : rom_o = 12'b110110001001; //2.792308
      780 : rom_o = 12'b110110110110; //2.828571
      781 : rom_o = 12'b110110110110; //2.828571
      782 : rom_o = 12'b110110110110; //2.828571
      783 : rom_o = 12'b110110110110; //2.828571
      784 : rom_o = 12'b110110110110; //2.828571
      785 : rom_o = 12'b110110110110; //2.828571
      786 : rom_o = 12'b110110110110; //2.828571
      787 : rom_o = 12'b110110110110; //2.828571
      788 : rom_o = 12'b110110110110; //2.828571
      789 : rom_o = 12'b110110110110; //2.828571
      790 : rom_o = 12'b110111100011; //2.864835
      791 : rom_o = 12'b110111100011; //2.864835
      792 : rom_o = 12'b110111100011; //2.864835
      793 : rom_o = 12'b110111100011; //2.864835
      794 : rom_o = 12'b110111100011; //2.864835
      795 : rom_o = 12'b110111100011; //2.864835
      796 : rom_o = 12'b110111100011; //2.864835
      797 : rom_o = 12'b110111100011; //2.864835
      798 : rom_o = 12'b110111100011; //2.864835
      799 : rom_o = 12'b110111100011; //2.864835
      800 : rom_o = 12'b111000010000; //2.901099
      801 : rom_o = 12'b111000010000; //2.901099
      802 : rom_o = 12'b111000010000; //2.901099
      803 : rom_o = 12'b111000010000; //2.901099
      804 : rom_o = 12'b111000010000; //2.901099
      805 : rom_o = 12'b111000010000; //2.901099
      806 : rom_o = 12'b111000010000; //2.901099
      807 : rom_o = 12'b111000010000; //2.901099
      808 : rom_o = 12'b111000010000; //2.901099
      809 : rom_o = 12'b111000010000; //2.901099
      810 : rom_o = 12'b111000111101; //2.937363
      811 : rom_o = 12'b111000111101; //2.937363
      812 : rom_o = 12'b111000111101; //2.937363
      813 : rom_o = 12'b111000111101; //2.937363
      814 : rom_o = 12'b111000111101; //2.937363
      815 : rom_o = 12'b111000111101; //2.937363
      816 : rom_o = 12'b111000111101; //2.937363
      817 : rom_o = 12'b111000111101; //2.937363
      818 : rom_o = 12'b111000111101; //2.937363
      819 : rom_o = 12'b111000111101; //2.937363
      820 : rom_o = 12'b111001101010; //2.973626
      821 : rom_o = 12'b111001101010; //2.973626
      822 : rom_o = 12'b111001101010; //2.973626
      823 : rom_o = 12'b111001101010; //2.973626
      824 : rom_o = 12'b111001101010; //2.973626
      825 : rom_o = 12'b111001101010; //2.973626
      826 : rom_o = 12'b111001101010; //2.973626
      827 : rom_o = 12'b111001101010; //2.973626
      828 : rom_o = 12'b111001101010; //2.973626
      829 : rom_o = 12'b111001101010; //2.973626
      830 : rom_o = 12'b111010010111; //3.009890
      831 : rom_o = 12'b111010010111; //3.009890
      832 : rom_o = 12'b111010010111; //3.009890
      833 : rom_o = 12'b111010010111; //3.009890
      834 : rom_o = 12'b111010010111; //3.009890
      835 : rom_o = 12'b111010010111; //3.009890
      836 : rom_o = 12'b111010010111; //3.009890
      837 : rom_o = 12'b111010010111; //3.009890
      838 : rom_o = 12'b111010010111; //3.009890
      839 : rom_o = 12'b111010010111; //3.009890
      840 : rom_o = 12'b111011000100; //3.046154
      841 : rom_o = 12'b111011000100; //3.046154
      842 : rom_o = 12'b111011000100; //3.046154
      843 : rom_o = 12'b111011000100; //3.046154
      844 : rom_o = 12'b111011000100; //3.046154
      845 : rom_o = 12'b111011000100; //3.046154
      846 : rom_o = 12'b111011000100; //3.046154
      847 : rom_o = 12'b111011000100; //3.046154
      848 : rom_o = 12'b111011000100; //3.046154
      849 : rom_o = 12'b111011000100; //3.046154
      850 : rom_o = 12'b111011110001; //3.082418
      851 : rom_o = 12'b111011110001; //3.082418
      852 : rom_o = 12'b111011110001; //3.082418
      853 : rom_o = 12'b111011110001; //3.082418
      854 : rom_o = 12'b111011110001; //3.082418
      855 : rom_o = 12'b111011110001; //3.082418
      856 : rom_o = 12'b111011110001; //3.082418
      857 : rom_o = 12'b111011110001; //3.082418
      858 : rom_o = 12'b111011110001; //3.082418
      859 : rom_o = 12'b111011110001; //3.082418
      860 : rom_o = 12'b111100011110; //3.118681
      861 : rom_o = 12'b111100011110; //3.118681
      862 : rom_o = 12'b111100011110; //3.118681
      863 : rom_o = 12'b111100011110; //3.118681
      864 : rom_o = 12'b111100011110; //3.118681
      865 : rom_o = 12'b111100011110; //3.118681
      866 : rom_o = 12'b111100011110; //3.118681
      867 : rom_o = 12'b111100011110; //3.118681
      868 : rom_o = 12'b111100011110; //3.118681
      869 : rom_o = 12'b111100011110; //3.118681
      870 : rom_o = 12'b111101001011; //3.154945
      871 : rom_o = 12'b111101001011; //3.154945
      872 : rom_o = 12'b111101001011; //3.154945
      873 : rom_o = 12'b111101001011; //3.154945
      874 : rom_o = 12'b111101001011; //3.154945
      875 : rom_o = 12'b111101001011; //3.154945
      876 : rom_o = 12'b111101001011; //3.154945
      877 : rom_o = 12'b111101001011; //3.154945
      878 : rom_o = 12'b111101001011; //3.154945
      879 : rom_o = 12'b111101001011; //3.154945
      880 : rom_o = 12'b111101111000; //3.191209
      881 : rom_o = 12'b111101111000; //3.191209
      882 : rom_o = 12'b111101111000; //3.191209
      883 : rom_o = 12'b111101111000; //3.191209
      884 : rom_o = 12'b111101111000; //3.191209
      885 : rom_o = 12'b111101111000; //3.191209
      886 : rom_o = 12'b111101111000; //3.191209
      887 : rom_o = 12'b111101111000; //3.191209
      888 : rom_o = 12'b111101111000; //3.191209
      889 : rom_o = 12'b111101111000; //3.191209
      890 : rom_o = 12'b111110100101; //3.227473
      891 : rom_o = 12'b111110100101; //3.227473
      892 : rom_o = 12'b111110100101; //3.227473
      893 : rom_o = 12'b111110100101; //3.227473
      894 : rom_o = 12'b111110100101; //3.227473
      895 : rom_o = 12'b111110100101; //3.227473
      896 : rom_o = 12'b111110100101; //3.227473
      897 : rom_o = 12'b111110100101; //3.227473
      898 : rom_o = 12'b111110100101; //3.227473
      899 : rom_o = 12'b111110100101; //3.227473
      900 : rom_o = 12'b111111010010; //3.263736
      901 : rom_o = 12'b111111010010; //3.263736
      902 : rom_o = 12'b111111010010; //3.263736
      903 : rom_o = 12'b111111010010; //3.263736
      904 : rom_o = 12'b111111010010; //3.263736
      905 : rom_o = 12'b111111010010; //3.263736
      906 : rom_o = 12'b111111010010; //3.263736
      907 : rom_o = 12'b111111010010; //3.263736
      908 : rom_o = 12'b111111010010; //3.263736
      909 : rom_o = 12'b111111010010; //3.263736
      910 : rom_o = 12'b111111111111; //3.300000
      911 : rom_o = 12'b111111111111; //3.300000
      912 : rom_o = 12'b111111111111; //3.300000
      913 : rom_o = 12'b111111111111; //3.300000
      914 : rom_o = 12'b111111111111; //3.300000
      915 : rom_o = 12'b111111111111; //3.300000
      916 : rom_o = 12'b111111111111; //3.300000
      917 : rom_o = 12'b111111111111; //3.300000
      918 : rom_o = 12'b111111111111; //3.300000
      919 : rom_o = 12'b111111111111; //3.300000
	  default: rom_o = 12'b000000000000;
	endcase
endmodule