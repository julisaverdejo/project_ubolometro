// Author: Julisa Verdejo Palacios
// Name: rom_volts.v
//
// Description: 


module rom_volts (
  input      [7:0] addr_i,
  output reg [11:0] rom_o
);

  always@(addr_i)  
    case(addr_i)
       0 : rom_o = 12'b000000000000; //0.000000
       1 : rom_o = 12'b000000101101; //0.036264
       2 : rom_o = 12'b000001011010; //0.072527
       3 : rom_o = 12'b000010000111; //0.108791
       4 : rom_o = 12'b000010110100; //0.145055
       5 : rom_o = 12'b000011100001; //0.181319
       6 : rom_o = 12'b000100001110; //0.217582
       7 : rom_o = 12'b000100111011; //0.253846
       8 : rom_o = 12'b000101101000; //0.290110
       9 : rom_o = 12'b000110010101; //0.326374
      10 : rom_o = 12'b000111000010; //0.362637
      11 : rom_o = 12'b000111101111; //0.398901
      12 : rom_o = 12'b001000011100; //0.435165
      13 : rom_o = 12'b001001001001; //0.471429
      14 : rom_o = 12'b001001110110; //0.507692
      15 : rom_o = 12'b001010100011; //0.543956
      16 : rom_o = 12'b001011010000; //0.580220
      17 : rom_o = 12'b001011111101; //0.616484
      18 : rom_o = 12'b001100101010; //0.652747
      19 : rom_o = 12'b001101010111; //0.689011
      20 : rom_o = 12'b001110000100; //0.725275
      21 : rom_o = 12'b001110110001; //0.761538
      22 : rom_o = 12'b001111011110; //0.797802
      23 : rom_o = 12'b010000001011; //0.834066
      24 : rom_o = 12'b010000111000; //0.870330
      25 : rom_o = 12'b010001100101; //0.906593
      26 : rom_o = 12'b010010010010; //0.942857
      27 : rom_o = 12'b010010111111; //0.979121
      28 : rom_o = 12'b010011101100; //1.015385
      29 : rom_o = 12'b010100011001; //1.051648
      30 : rom_o = 12'b010101000110; //1.087912
      31 : rom_o = 12'b010101110011; //1.124176
      32 : rom_o = 12'b010110100000; //1.160440
      33 : rom_o = 12'b010111001101; //1.196703
      34 : rom_o = 12'b010111111010; //1.232967
      35 : rom_o = 12'b011000100111; //1.269231
      36 : rom_o = 12'b011001010100; //1.305495
      37 : rom_o = 12'b011010000001; //1.341758
      38 : rom_o = 12'b011010101110; //1.378022
      39 : rom_o = 12'b011011011011; //1.414286
      40 : rom_o = 12'b011100001000; //1.450549
      41 : rom_o = 12'b011100110101; //1.486813
      42 : rom_o = 12'b011101100010; //1.523077
      43 : rom_o = 12'b011110001111; //1.559341
      44 : rom_o = 12'b011110111100; //1.595604
      45 : rom_o = 12'b011111101001; //1.631868
      46 : rom_o = 12'b100000010110; //1.668132
      47 : rom_o = 12'b100001000011; //1.704396
      48 : rom_o = 12'b100001110000; //1.740659
      49 : rom_o = 12'b100010011101; //1.776923
      50 : rom_o = 12'b100011001010; //1.813187
      51 : rom_o = 12'b100011110111; //1.849451
      52 : rom_o = 12'b100100100100; //1.885714
      53 : rom_o = 12'b100101010001; //1.921978
      54 : rom_o = 12'b100101111110; //1.958242
      55 : rom_o = 12'b100110101011; //1.994505
      56 : rom_o = 12'b100111011000; //2.030769
      57 : rom_o = 12'b101000000101; //2.067033
      58 : rom_o = 12'b101000110010; //2.103297
      59 : rom_o = 12'b101001011111; //2.139560
      60 : rom_o = 12'b101010001100; //2.175824
      61 : rom_o = 12'b101010111001; //2.212088
      62 : rom_o = 12'b101011100110; //2.248352
      63 : rom_o = 12'b101100010011; //2.284615
      64 : rom_o = 12'b101101000000; //2.320879
      65 : rom_o = 12'b101101101101; //2.357143
      66 : rom_o = 12'b101110011010; //2.393407
      67 : rom_o = 12'b101111000111; //2.429670
      68 : rom_o = 12'b101111110100; //2.465934
      69 : rom_o = 12'b110000100001; //2.502198
      70 : rom_o = 12'b110001001110; //2.538462
      71 : rom_o = 12'b110001111011; //2.574725
      72 : rom_o = 12'b110010101000; //2.610989
      73 : rom_o = 12'b110011010101; //2.647253
      74 : rom_o = 12'b110100000010; //2.683516
      75 : rom_o = 12'b110100101111; //2.719780
      76 : rom_o = 12'b110101011100; //2.756044
      77 : rom_o = 12'b110110001001; //2.792308
      78 : rom_o = 12'b110110110110; //2.828571
      79 : rom_o = 12'b110111100011; //2.864835
      80 : rom_o = 12'b111000010000; //2.901099
      81 : rom_o = 12'b111000111101; //2.937363
      82 : rom_o = 12'b111001101010; //2.973626
      83 : rom_o = 12'b111010010111; //3.009890
      84 : rom_o = 12'b111011000100; //3.046154
      85 : rom_o = 12'b111011110001; //3.082418
      86 : rom_o = 12'b111100011110; //3.118681
      87 : rom_o = 12'b111101001011; //3.154945
      88 : rom_o = 12'b111101111000; //3.191209
      89 : rom_o = 12'b111110100101; //3.227473
      90 : rom_o = 12'b111111010010; //3.263736
      91 : rom_o = 12'b111111111111; //3.300000	  
	  
	  default: rom_o = 12'b000000000000;
	endcase
endmodule